library library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity alu is
    port (
        s0, s1, s2, i0, i1, j0, j1 : in std_logic;
        k0, k1, c_out : out std_logic
    );
end entity alu;

architecture struc of alu is
    
begin
    
    
    
end architecture struc;